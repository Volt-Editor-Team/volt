module list

pub struct ListCursor {
}
