module ui

// import core.controller as ctl

pub enum Ui {
	tui
	gui
}

// pub fn initialize(ui_design Ui) {
// 	match ui_design {
// 		.tui {
// 			return
// 		}
// 	}
// }
