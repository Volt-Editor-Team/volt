module cursor
