module core

pub const default_tabsize = 4
