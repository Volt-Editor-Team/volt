module tui

// import core.controller
// import term

fn draw_changes(x voidptr) {
	// width, height := term.get_terminal_size()

	// // get app pointer, terminal size, and clear to prep for updates
	// mut tui_app := get_tui(x)
	// mut ctx := tui_app.tui
	// mut app := controller.get_app(tui_app.core)

	// // relavent info for rendering
	// mut view := &app.viewport
	// mut buf := app.buffers[app.active_buffer]
}
