module gap

fn test_delete() {
	mut buf := GapBuffer.new(GapBuffer{})
	assert buf.to_string() == ''
	assert buf.debug_string() == '[gap:0]'
	buf.insert(2, '2345678')
	assert buf.to_string() == '2345678'
	assert buf.debug_string() == '2345678[gap:7]'
	buf.delete(2, 3)
	assert buf.to_string() == '2378'
	assert buf.debug_string() == '23[gap:10]78'
	buf.delete(0, 1)
	assert buf.to_string() == '378'
	assert buf.debug_string() == '[gap:11]378'
}
