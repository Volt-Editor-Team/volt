module tui

import core.controller as ctl
import term.ui as t

pub fn get_tui(x voidptr) &TuiApp {
	return unsafe { &TuiApp(x) }
}

pub struct TuiApp {
pub mut:
	core  voidptr
	tui   &TuiContext = unsafe { nil }
	theme TuiTheme
}

type TuiContext = t.Context

pub fn TuiApp.new(core voidptr) &TuiApp {
	mut tui_app := &TuiApp{}
	tui_app.initialize_tui(core)

	return tui_app
}

pub fn (mut tui_app TuiApp) initialize_tui(core voidptr) {
	tui_app.core = core
	app := ctl.get_app(core)
	tui_app.theme = TuiTheme.new(app.theme)
	tui_app.tui = t.init(
		init_fn:        full_redraw
		user_data:      tui_app
		event_fn:       event_wrapper
		frame_fn:       full_redraw
		capture_events: true
		hide_cursor:    true
		frame_rate:     30
	)
}

pub fn event_wrapper(e &t.Event, x voidptr) {
	tui_app := get_tui(x)
	event_type := convert_event_type(e.typ)
	key_code := convert_key_code(e.code)
	modifier := convert_modifier(e.modifiers)
	input := ctl.UserInput{
		mod:  modifier
		e:    event_type
		code: key_code
	}

	ctl.event_loop(input, tui_app.core)
}
