module viewport

pub fn (mut view Viewport) update_visual_wraps(x int) {
	view.visual_wraps = x
}
