module viewport

pub struct Viewport {
pub mut:
	row_offset int
	col_offset int
pub:
	height int
	width  int
	margin int
}
