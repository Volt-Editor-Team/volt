module rope

import gap

fn test_iterator() {
}
