module viewport
