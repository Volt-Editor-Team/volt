module controller

import fs
import os
import util
import math
import time

pub fn handle_normal_mode_event(x voidptr, mod Modifier, event EventType, key KeyCode) {
	mut app := get_app(x)
	mut buf := &app.buffers[app.active_buffer]
	mut view := &app.viewport
	// global normal mode
	if event == .key_down {
		if buf.cmd.command.len > 0 {
			buf.cmd.command = ''
		}
		match key {
			.f {
				buf.change_mode(.search, true)
			}
			.space {
				buf.change_mode(.menu, true)
			}
			.g {
				buf.change_mode(.goto, true)
			}
			.i {
				buf.change_mode(.insert, false)
			}
			.colon {
				buf.change_mode(.command, false)
			}
			else {}
		}
	}

	// specific to persistant mode
	if buf.p_mode == .default || buf.p_mode == .directory {
		if event == .key_down {
			match key {
				.d {
					// currently just deletes one character
					// will need to be changed when selections are supported
					buf.delete(view.cursor.flat_index, 1)
					updated_line := buf.buffer.line_at(view.cursor.y).clone()
					view.visible_lines[view.cursor.y - view.row_offset] = updated_line
				}
				.l, .right {
					prev_y := view.cursor.y
					view.cursor.move_right_buffer(view.visible_lines, view.row_offset,
						view.tabsize)
					view.cursor.update_desired_col(app.viewport.width)

					if view.cursor.y != prev_y {
						view.update_offset(view.cursor.y, buf.buffer)
					}
				}
				.h, .left {
					prev_y := view.cursor.y
					view.cursor.move_left_buffer(view.visible_lines, view.row_offset,
						view.tabsize)
					view.cursor.update_desired_col(app.viewport.width)
					if view.cursor.y != prev_y {
						view.update_offset(view.cursor.y, buf.buffer)
						// buf.update_offset(app.viewport.visual_wraps, app.viewport.height,
						// 	app.viewport.margin, app.viewport.row_offset)
					}
				}
				.j, .down {
					line := view.visible_lines[view.cursor.y - view.row_offset]

					// total wraps in the current line
					mut total_wraps := 0
					if line.len != 0 {
						total_wraps = util.char_count_expanded_tabs(line, view.tabsize) / app.viewport.width
					}

					// current wrap index
					cur_wrap := view.cursor.visual_x / app.viewport.width

					if cur_wrap < total_wraps {
						mut perfect_index := util.expand_tabs_to(line#[..view.cursor.x +
							app.viewport.width - 1], view.cursor.x + app.viewport.width - 1,
							view.tabsize)
						if view.cursor.x + app.viewport.width - 1 <= line.len {
							perfect_index++
						}
						view.cursor.move_to_x(line, perfect_index, view.tabsize)
					} else {
						view.cursor.move_down_buffer(view.visible_lines, view.row_offset,
							view.tabsize)
					}

					// update viewport offset
					view.update_offset(view.cursor.y, buf.buffer)
				}
				.k, .up {
					relative_y := view.cursor.y - view.row_offset
					cur_wrap := util.char_count_expanded_tabs(view.visible_lines[relative_y]#[..view.cursor.x],
						view.tabsize) / app.viewport.width
					if cur_wrap == 0 {
						// line above is NOT the first line
						if view.cursor.y - 1 > 0 {
							line := view.visible_lines[relative_y - 1]

							mut total_wraps := 0
							if line.len != 0 {
								total_wraps = util.char_count_expanded_tabs(line, view.tabsize) / app.viewport.width
							}
							if total_wraps > 0 {
								view.cursor.move_up_buffer(view.visible_lines, view.row_offset,
									view.tabsize)
								mut index := total_wraps * app.viewport.width + view.cursor.x
								perfect_index := util.expand_tabs_to(line#[..index - 1],
									index - 1, view.tabsize)
								view.cursor.move_to_x(buf.cur_line, perfect_index, view.tabsize)
							} else {
								view.cursor.move_up_buffer(view.visible_lines, view.row_offset,
									view.tabsize)
							}
						} else {
							view.cursor.move_up_buffer(view.visible_lines, view.row_offset,
								view.tabsize)
						}
					} else {
						line := view.visible_lines[relative_y]
						index := math.max(cur_wrap * app.viewport.width + view.cursor.desired_col,
							view.cursor.x)
						next_index := util.expand_tabs_to(line#[..index - app.viewport.width - 1],
							index - app.viewport.width - 1, view.tabsize)
						view.cursor.move_to_x(buf.cur_line, math.min(next_index, view.cursor.desired_col),
							view.tabsize)
					}

					// update offset
					view.update_offset(view.cursor.y, buf.buffer)
				}
				else {}
			}
		}
	}
	match buf.p_mode {
		.directory {
			match mod {
				.none {
					match key {
						.enter {
							path := buf.buffer.line_at(view.cursor.y).string()
							app.add_new_buffer(
								name: os.file_name(path)
								path: buf.path + path
								// tabsize: view.tabsize
								type:   .gap
								mode:   .normal
								p_mode: .default
							)
						}
						.tab {
							path := buf.buffer.line_at(view.cursor.y).string()

							if fs.is_dir(buf.path + path) {
								parent_dir, paths := fs.get_paths_from_dir(buf.path, path)
								buf.path = parent_dir
								replacement_runes := [][]rune{len: paths.len, init: paths[index].runes()}
								buf.buffer.replace_with_temp(replacement_runes)

								view.cursor.x = 0
								view.cursor.y = 0
								view.cursor.flat_index = 0
							}
						}
						.backspace {
							parent_dir, paths := fs.get_paths_from_parent_dir(buf.path)
							buf.path = parent_dir
							replacement_runes := [][]rune{len: paths.len, init: paths[index].runes()}
							buf.buffer.replace_with_temp(replacement_runes)

							view.cursor.x = 0
							view.cursor.y = 0
							view.cursor.flat_index = 0
						}
						else {}
					}
				}
				else {}
			}
		}
		.fuzzy {
			match mod {
				.none {
					match key {
						.escape {
							// restore settings
							buf.p_mode = buf.temp_mode
							buf.change_mode(.normal, false)
							view.update_offset(view.cursor.y, buf.buffer)
							view.fill_visible_lines(buf.buffer)

							// delete temp stuff
							// buf.temp_label = ''
							// buf.temp_data.clear()
							buf.clear_all_temp_data()
							buf.file_ch.close()
						}
						.j, .down {
							if buf.temp_cursor.y < buf.temp_data.len - 1 {
								buf.temp_cursor.y++
								view.update_offset_for_temp(buf.temp_cursor.y)
							}
						}
						.k, .up {
							if buf.temp_cursor.y > 0 {
								buf.temp_cursor.y--
								view.update_offset_for_temp(buf.temp_cursor.y)
							}
						}
						// for switch fuzzy search directory
						.tab {
							if buf.temp_data.len > 0 {
								file := buf.temp_data[buf.temp_cursor.y].string()

								path := buf.temp_path + os.path_separator + file

								if os.is_dir(path) {
									buf.temp_path = path
									// delete temp stuff
									buf.temp_label = ''
									buf.temp_data.clear()
									buf.file_ch.close()
									buf.p_mode = buf.temp_mode
									buf.temp_fuzzy_type = .dir
									// reset and open fuzzy
									buf.open_fuzzy_find(buf.temp_path, .directory)
									time.sleep(80 * time.millisecond)
									buf.temp_cursor.y = math.min(buf.temp_data.len - 1,
										buf.temp_cursor.y)
									view.update_offset_for_temp(buf.temp_cursor.y)
								}
							}
						}
						.backtick {
							if buf.temp_fuzzy_type == .dir {
								buf.temp_label = ''
								buf.temp_data.clear()
								buf.file_ch.close()
								buf.p_mode = buf.temp_mode
								buf.temp_fuzzy_type = .file
								// reset and open fuzzy
								buf.open_fuzzy_find(buf.temp_path, .file)
								time.sleep(80 * time.millisecond)
								buf.temp_cursor.y = math.min(buf.temp_data.len - 1, buf.temp_cursor.y)
								view.update_offset_for_temp(buf.temp_cursor.y)
							} else if buf.temp_fuzzy_type == .file {
								buf.temp_label = ''
								buf.temp_data.clear()
								buf.file_ch.close()
								buf.p_mode = buf.temp_mode
								buf.temp_fuzzy_type = .dir
								// reset and open fuzzy
								buf.open_fuzzy_find(buf.temp_path, .directory)
								time.sleep(80 * time.millisecond)
								buf.temp_cursor.y = math.min(buf.temp_data.len - 1, buf.temp_cursor.y)
								view.update_offset_for_temp(buf.temp_cursor.y)
							}
						}
						.o {
							if buf.temp_data.len > 0 {
								file := buf.temp_data[buf.temp_cursor.y].string()

								path := buf.temp_path + os.path_separator + file

								if os.is_dir(path) {
									buf.temp_path = path
									// delete temp stuff
									buf.temp_label = ''
									buf.temp_int = 0
									buf.temp_data.clear()
									buf.file_ch.close()
									// reset and open fuzzy
									buf.p_mode = buf.temp_mode
									buf.temp_fuzzy_type = .file
									buf.open_fuzzy_find(buf.temp_path, .file)
									time.sleep(80 * time.millisecond)
									buf.temp_cursor.y = math.min(buf.temp_data.len - 1,
										buf.temp_cursor.y)
									view.update_offset_for_temp(buf.temp_cursor.y)
								}
							}
						}
						.comma {
							if buf.temp_data.len > 0 {
								if buf.temp_cursor.y < 0
									|| buf.temp_cursor.y > buf.temp_data.len - 1 {
									buf.temp_cursor.y = math.min(buf.temp_data.len - 1,
										buf.temp_cursor.y)
								}
								file := buf.temp_data[buf.temp_cursor.y].string()
								mut path := buf.temp_path + os.path_separator + file

								if os.is_file(path) {
									if buf.temp_list.contains(path) {
										mut index := 0
										for p in buf.temp_list {
											if p == path {
												break
											}
											index++
										}
										buf.temp_list.delete(index)
									} else {
										buf.temp_list << path
									}
									buf.temp_label = ''
								}
							}
						}
						.enter {
							if buf.temp_data.len > 0 {
								file := buf.temp_data[buf.temp_cursor.y].string()

								// buf.path = buf.temp_path
								buf.p_mode = buf.temp_mode
								buf.mode = .normal
								// buf.logical_cursor = buf.temp_cursor
								view.update_offset(view.cursor.y, buf.buffer)
								view.existing_cursors[app.active_buffer] = view.cursor
								view.existing_offsets[app.active_buffer] = view.row_offset
								buf.file_ch.close()

								// delete temp stuff
								mut path := buf.temp_path + os.path_separator + file

								if os.is_dir(path) {
									dir_path := path + os.path_separator
									for mut buffer in app.buffers {
										full_path := app.working_dir + os.path_separator +
											buffer.path
										if full_path.starts_with(dir_path) {
											buffer.path = full_path.replace(dir_path,
												'')
										} else {
											buffer.path = full_path
										}
									}
									os.chdir(path) or { return }
									app.working_dir = path
								} else {
									buf.temp_list << path
									// if buf.temp_list.len == 0 {
									// 	buf.temp_list << path
									// }
								}
								file_list := buf.temp_list.clone()
								// tabsize := view.tabsize

								for i, paths in file_list {
									if i == 0 {
										app.add_new_buffer(
											name: os.file_name(paths)
											path: paths
											// tabsize: tabsize
											type:   .gap
											mode:   .normal
											p_mode: .default
										)
									} else {
										app.append_new_buffer(
											name: os.file_name(paths)
											path: paths
											// tabsize: tabsize
											type:   .gap
											mode:   .normal
											p_mode: .default
										)
									}
								}
								app.active_buffer = app.buffers.len - 1
								view.row_offset = if view.existing_offsets.keys().contains(app.active_buffer) {
									view.existing_offsets[app.active_buffer]
								} else {
									0
								}
								if view.existing_cursors.keys().contains(app.active_buffer) {
									view.cursor = view.existing_cursors[app.active_buffer]
								} else {
									view.cursor.x = 0
									view.cursor.y = 0
									view.cursor.flat_index = 0
									view.cursor.visual_x = 0
									view.cursor.desired_col = 0
								}

								view.fill_visible_lines(app.buffers[app.active_buffer].buffer)
								// view.fill_visible_lines(buf.buffer)
								buf.temp_list.clear()
								buf.temp_label = ''
								buf.temp_int = 0
								buf.temp_data.clear()
								buf.menu_state = false
							}
						}
						else {}
					}
				}
				.shift {
					match key {
						// for switch fuzzy search directory
						.tab {
							buf.temp_path = os.dir(buf.temp_path)
							if os.is_dir(buf.temp_path) {
								// delete temp stuff
								buf.temp_label = ''
								buf.temp_int = 0
								buf.temp_data.clear()
								buf.file_ch.close()
								buf.p_mode = buf.temp_mode
								buf.temp_fuzzy_type = .dir
								// reset and open fuzzy
								buf.open_fuzzy_find(buf.temp_path, .directory)
								// buf.temp_cursor.y = 0
								time.sleep(80 * time.millisecond)
								buf.temp_cursor.y = math.min(buf.temp_data.len - 1, buf.temp_cursor.y)
								view.update_offset_for_temp(buf.temp_cursor.y)
							}
						}
						else {}
					}
				}
				else {}
			}
		}
		else {}
	}
}
