module util

import term.ui as tui

pub const neutral_grey = tui.Color{
	r: 38
	g: 50
	b: 56
}

pub const teal = tui.Color{
	r: 0
	g: 150
	b: 136
}

pub const amber = tui.Color{
	r: 255
	g: 171
	b: 64
}

pub const purple = tui.Color{
	r: 156
	g: 36
	b: 176
}

pub const deep_indigo = tui.Color{
	r: 63
	g: 81
	b: 181
}
